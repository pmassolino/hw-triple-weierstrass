----------------------------------------------------------------------------------
-- Engineer: Pedro Maat C. Massolino
-- 
-- Create Date:    11/11/2016
-- Design Name:    controller_small_montgomery_processor_3
-- Module Name:    controller_small_montgomery_processor_3
-- Project Name:   Montgomery processor
-- Target Devices: Any
-- Tool versions:  Microsemi Libero 11.7
--
-- Description: 
--
-- This is the state machine that controls the Montgomery processor unit.
-- It can handle all these instructions:
-- 
-- Multiplication Instruction (000)
-- Performs the Montgomery multiplication of two values.
-- It has to be performed on two variables that can be equal.
-- But the output has to be different. Also, the variable 0 is always the prime.
-- a*b -> p
-- 'a' can be equal to 'b', but 'p' has to be different than both of them.
--
-- Addition Instruction (001)
-- Performs the addition of two numbers without reducing the modulo of the prime.
-- This can be performed by the same variable as input.
-- However variable 'b' has to be the same as the output variable 'p'.
-- b + a -> p
--
-- Subtraction Normalized Instruction (010)
-- Performs the subtraction of two values and add the prime multiplied by a constant.
-- This addition of the prime guarantee the output is not negative.
-- This can be performed by the same variable as input.
-- However variable 'b' has to be the same as the output variable 'p'.
-- b - a -> p
-- Also only variable in 'a' can be negative.
--
-- Subtraction Instruction (011)
-- Performs subtraction of two values without reducing or normalizing.
-- The rule is the same as the subtraction with normalization. 
-- b - a -> p
--
--
-- Do nothing (111)
--
--
-- Dependencies:
-- VHDL-93
--
-- 
-- Revision: 
-- Revision 1.0
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity controller_small_montgomery_processor_3 is
    Port(
        clk : in STD_LOGIC;
        rst : in STD_LOGIC;
        start : in STD_LOGIC;
        counters_limit : in STD_LOGIC;
        instruction : in STD_LOGIC_VECTOR(2 downto 0);
        mem_write_enable_new_value : out STD_LOGIC;
        reg_processor_free_d : out STD_LOGIC;
        reg_operands_size_ce : out STD_LOGIC;
        reg_variables_ce : out STD_LOGIC;
        counter_a_j_ce : out STD_LOGIC;
        counter_a_j_rst : out STD_LOGIC;
        counter_b_i_ce : out STD_LOGIC;
        counter_b_i_rst : out STD_LOGIC;
        address_n_ce : out STD_LOGIC;
        address_n_load : out STD_LOGIC;
        address_n_rst : out STD_LOGIC;
        address_new_p_ce : out STD_LOGIC;
        address_new_p_rst : out STD_LOGIC;
        dsp1_a_en : out STD_LOGIC;
        dsp1_a_rst : out STD_LOGIC;
        reg_b_ce : out STD_LOGIC;
        reg_b_rst : out STD_LOGIC;
        dsp1_c_en : out STD_LOGIC;
        dsp1_c_rst : out STD_LOGIC;
        dsp1_add_sub_mode : out STD_LOGIC;
        dsp1_reg_add_sub_mode_ce : out STD_LOGIC;
        dsp1_accumulation_mode : out STD_LOGIC;
        dsp1_reg_accumulation_mode_ce : out STD_LOGIC;
        dsp1_external_carry_in_mode : out STD_LOGIC;
        dsp1_reg_external_carry_in_mode_ce : out STD_LOGIC;
        dsp1_arshift_mode : out STD_LOGIC;
        dsp1_reg_arshift_mode_ce : out STD_LOGIC;
        dsp1_p_en : out STD_LOGIC;
        dsp1_p_rst : out STD_LOGIC;
        reg_m_ce : out STD_LOGIC;
        reg_m_rst : out STD_LOGIC;
        dsp2_b_en : out STD_LOGIC;
        dsp2_b_rst : out STD_LOGIC;
        dsp2_c_en : out STD_LOGIC;
        dsp2_c_rst : out STD_LOGIC;
        dsp2_add_sub_mode : out STD_LOGIC;
        dsp2_reg_add_sub_mode_ce : out STD_LOGIC;
        dsp2_accumulation_mode : out STD_LOGIC;
        dsp2_reg_accumulation_mode_ce : out STD_LOGIC;
        dsp2_external_carry_in_mode : out STD_LOGIC;
        dsp2_reg_external_carry_in_mode_ce : out STD_LOGIC;
        dsp2_arshift_mode : out STD_LOGIC;
        dsp2_reg_arshift_mode_ce : out STD_LOGIC;
        dsp2_p_en : out STD_LOGIC;
        dsp2_p_rst : out STD_LOGIC;
        sel_load_b_i : out STD_LOGIC;
        sel_value_m : out STD_LOGIC;
        sel_compare_counter_b_i : out STD_LOGIC
    );
end controller_small_montgomery_processor_3;

architecture Behavioral of controller_small_montgomery_processor_3 is

component register_rst_nbits
    Generic (size : integer);
    Port (
        d : in STD_LOGIC_VECTOR ((size - 1) downto 0);
        clk : in STD_LOGIC;
        ce : in STD_LOGIC;
        rst : in STD_LOGIC;
        rst_value : in STD_LOGIC_VECTOR ((size - 1) downto 0);
        q : out  STD_LOGIC_VECTOR ((size - 1) downto 0)
    );
end component;

type State is (reset, decode_instruction,
-- Multiplication Instruction States
begin_montgomery_multiplication,
begin_reset_counters_montgomery_multiplication, load_registers_1_first_iteration_montgomery_multiplication, load_registers_2_first_iteration_montgomery_multiplication, prepare_compute_m_1_first_iteration_montgomery_multiplication, prepare_compute_m_2_first_iteration_montgomery_multiplication, compute_m_first_iteration_montgomery_multiplication, prepare_compute_1_first_iteration_montgomery_multiplication, prepare_compute_2_first_iteration_montgomery_multiplication, prepare_compute_3_first_iteration_montgomery_multiplication, compute_first_iteration_montgomery_multiplication, last_compute_1_first_iteration_montgomery_multiplication, last_compute_2_first_iteration_montgomery_multiplication, last_compute_3_first_iteration_montgomery_multiplication,
last_compute_2_remaining_iterations_montgomery_multiplication, last_compute_3_remaining_iterations_montgomery_multiplication, last_compute_4_remaining_iterations_montgomery_multiplication, prepare_compute_m_1_remaining_iterations_montgomery_multiplication, prepare_compute_m_2_remaining_iterations_montgomery_multiplication, compute_m_remaining_iterations_montgomery_multiplication, prepare_compute_1_remaining_iterations_montgomery_multiplication, prepare_compute_2_remaining_iterations_montgomery_multiplication, prepare_compute_3_remaining_iterations_montgomery_multiplication, compute_remaining_iterations_montgomery_multiplication, last_compute_1_remaining_iterations_montgomery_multiplication,
last_compute_2_last_iterations_montgomery_multiplication, last_compute_3_last_iteration_montgomery_multiplication, last_compute_4_last_iteration_montgomery_multiplication, last_compute_5_last_iteration_montgomery_multiplication, last_compute_6_last_iteration_montgomery_multiplication, last_compute_7_last_iteration_montgomery_multiplication,  
finished_montgomery_multiplication,
-- Addition/Subtraction Instruction States
begin_montgomery_addition_subtraction_no_reduction,
begin_reset_counters_montgomery_addition_subtraction_no_reduction, prepare_compute_1_montgomery_addition_subtraction_no_reduction, prepare_compute_2_montgomery_addition_subtraction_no_reduction, prepare_compute_3_montgomery_addition_subtraction_no_reduction, prepare_compute_4_montgomery_addition_subtraction_no_reduction, compute_montgomery_addition_subtraction_no_reduction, last_compute_1_montgomery_addition_subtraction_no_reduction, last_compute_2_montgomery_addition_subtraction_no_reduction, last_compute_3_montgomery_addition_subtraction_no_reduction, last_compute_4_montgomery_addition_subtraction_no_reduction, last_compute_5_montgomery_addition_subtraction_no_reduction, last_compute_6_montgomery_addition_subtraction_no_reduction,
finished_montgomery_addition_subtraction_no_reduction
); 
signal actual_state, next_state : State;


signal reg_addition_subtraction_mode_d : STD_LOGIC_VECTOR(1 downto 0);
signal reg_addition_subtraction_mode_ce : STD_LOGIC;
constant reg_addition_subtraction_mode_rst_value : STD_LOGIC_VECTOR(1 downto 0) := "11";
signal reg_addition_subtraction_mode_q : STD_LOGIC_VECTOR(1 downto 0);

begin

Clock : process (clk)
begin
    if (rising_edge(clk)) then
        if(rst = '0') then
            actual_state <= reset;
        else
            actual_state <= next_state;
        end if;
    else
        null;
    end if;
end process;

Output : process (actual_state, start, instruction, reg_addition_subtraction_mode_q)
begin
    mem_write_enable_new_value <= '0';
    reg_processor_free_d <= '0';
    reg_addition_subtraction_mode_d <= "11";
    reg_addition_subtraction_mode_ce <= '0';
    reg_operands_size_ce <= '0';
    reg_variables_ce <= '0';
    counter_a_j_ce <= '0';
    counter_a_j_rst <= '1';
    counter_b_i_ce <= '0';
    counter_b_i_rst <= '1';
    address_n_ce <= '0';
    address_n_load <= '0';
    address_n_rst <= '1';
    address_new_p_ce <= '0';
    address_new_p_rst <= '1';
    dsp1_a_en <= '0';
    dsp1_a_rst <= '1';
    reg_b_ce <= '0';
    reg_b_rst <= '1';
    dsp1_c_en <= '0';
    dsp1_c_rst <= '1';
    dsp1_add_sub_mode <= '0';
    dsp1_reg_add_sub_mode_ce <= '0';
    dsp1_accumulation_mode <= '0';
    dsp1_reg_accumulation_mode_ce <= '0';
    dsp1_external_carry_in_mode <= '0';
    dsp1_reg_external_carry_in_mode_ce <= '0';
    dsp1_arshift_mode <= '0';
    dsp1_reg_arshift_mode_ce <= '0';
    dsp1_p_en <= '0';
    dsp1_p_rst <= '1';
    reg_m_ce <= '0';
    reg_m_rst <= '1';
    dsp2_b_en <= '0';
    dsp2_b_rst <= '1';
    dsp2_c_en <= '0';
    dsp2_c_rst <= '1';
    dsp2_add_sub_mode <= '0';
    dsp2_reg_add_sub_mode_ce <= '0';
    dsp2_accumulation_mode <= '0';
    dsp2_reg_accumulation_mode_ce <= '0';
    dsp2_external_carry_in_mode <= '0';
    dsp2_reg_external_carry_in_mode_ce <= '0';
    dsp2_arshift_mode <= '0';
    dsp2_reg_arshift_mode_ce <= '0';
    dsp2_p_en <= '0';
    dsp2_p_rst <= '1';
    sel_load_b_i <= '0';
    sel_value_m <= '0';
    sel_compare_counter_b_i <= '0';
    case (actual_state) is
        when reset =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';            
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '0';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '0';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '0';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '0';
            reg_b_ce <= '0';
            reg_b_rst <= '0';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '0';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '1';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '1';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '1';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '1';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '0';
            reg_m_ce <= '0';
            reg_m_rst <= '0';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '0';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '0';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '1';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '1';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '1';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '1';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '0';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when decode_instruction =>
            if(start = '0' or instruction = "111") then
                reg_operands_size_ce <= '0';
                reg_variables_ce <= '0';
            else
                reg_operands_size_ce <= '1';
                reg_variables_ce <= '1';
            end if;
            if(instruction = "001") then
                reg_addition_subtraction_mode_d <= "10";
                reg_addition_subtraction_mode_ce <= '1';
            elsif(instruction = "010") then
                reg_addition_subtraction_mode_d <= "01";
                reg_addition_subtraction_mode_ce <= '1';
            elsif(instruction = "011") then
                reg_addition_subtraction_mode_d <= "00";
                reg_addition_subtraction_mode_ce <= '1';
            else
                reg_addition_subtraction_mode_d <= "11";
                reg_addition_subtraction_mode_ce <= '1';
            end if;
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '1';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when begin_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '0';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '0';
            address_n_ce <= '1';
            address_n_load <= '1';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '0';
            reg_b_ce <= '0';
            reg_b_rst <= '0';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '0';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '1';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '1';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '1';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '1';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '0';
            reg_m_ce <= '0';
            reg_m_rst <= '0';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '0';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '0';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '1';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '1';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '1';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '1';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '0';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when begin_reset_counters_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '1';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when load_registers_1_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '1';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when load_registers_2_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '0';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '1';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '1';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '1';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '1';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_m_1_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_m_2_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '0';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '1';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '0';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '1';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '1';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '1';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '1';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when compute_m_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '1';
            dsp1_accumulation_mode <= '1';
            dsp1_reg_accumulation_mode_ce <= '1';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '1';
            dsp1_arshift_mode <= '1';
            dsp1_reg_arshift_mode_ce <= '1';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_1_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '1';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '1';
            dsp2_accumulation_mode <= '1';
            dsp2_reg_accumulation_mode_ce <= '1';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '1';
            dsp2_arshift_mode <= '1';
            dsp2_reg_arshift_mode_ce <= '1';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '0';
            sel_load_b_i <= '0';
            sel_value_m <= '1';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_2_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_3_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0'; 
        when compute_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';         
        when last_compute_1_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '0';
            counter_b_i_ce <= '1';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_2_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '0';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '1';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_3_first_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '0';
            reg_b_ce <= '1';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_4_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '1';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '1';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '1';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '1';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '0';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_m_1_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_m_2_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '0';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '1';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '0';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '1';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '1';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '1';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '1';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when compute_m_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '1';
            dsp1_accumulation_mode <= '1';
            dsp1_reg_accumulation_mode_ce <= '1';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '1';
            dsp1_arshift_mode <= '1';
            dsp1_reg_arshift_mode_ce <= '1';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_1_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '1';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '1';
            dsp2_accumulation_mode <= '1';
            dsp2_reg_accumulation_mode_ce <= '1';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '1';
            dsp2_arshift_mode <= '1';
            dsp2_reg_arshift_mode_ce <= '1';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '0';
            sel_load_b_i <= '0';
            sel_value_m <= '1';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_2_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_3_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when compute_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_1_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '1';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '1';
        when last_compute_2_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '0';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '0';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '1';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_3_remaining_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '1';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '0';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_2_last_iterations_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '0';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '0';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '1';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_3_last_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '0';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_4_last_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '0';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_5_last_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_6_last_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_7_last_iteration_montgomery_multiplication =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '1';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when finished_montgomery_multiplication =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '1';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '0';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '0';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '0';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '0';
            reg_b_ce <= '0';
            reg_b_rst <= '0';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '0';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '0';
            reg_m_ce <= '1';
            reg_m_rst <= '0';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '0';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '0';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '0';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when begin_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '0';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '0';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '0';
            reg_b_ce <= '0';
            reg_b_rst <= '0';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '0';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '0';
            reg_m_ce <= '0';
            reg_m_rst <= '0';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '0';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '0';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '0';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when begin_reset_counters_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_1_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '0';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            if(reg_addition_subtraction_mode_q(1) = '0') then
                dsp1_add_sub_mode <= '1';
            else
                dsp1_add_sub_mode <= '0';
            end if;
            dsp1_reg_add_sub_mode_ce <= '1';
            dsp1_accumulation_mode <= '1';
            dsp1_reg_accumulation_mode_ce <= '1';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '1';
            dsp1_arshift_mode <= '1';
            dsp1_reg_arshift_mode_ce <= '1';            
            dsp1_p_en <= '1';
            dsp1_p_rst <= '0';
            reg_m_ce <= '0';
            reg_m_rst <= '0';
            dsp2_b_en <= '1';
            dsp2_b_rst <= '0';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_2_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_3_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            if(reg_addition_subtraction_mode_q(0) = '0') then
                dsp2_b_en <= '0';
            else
                dsp2_b_en <= '1';
            end if;
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            if(reg_addition_subtraction_mode_q(1) = '0') then
                dsp2_accumulation_mode <= '1';
                dsp2_arshift_mode <= '1';
            else
                dsp2_accumulation_mode <= '0';
                dsp2_arshift_mode <= '0';
            end if;
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '1';
            dsp2_reg_accumulation_mode_ce <= '1';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '1';
            dsp2_reg_arshift_mode_ce <= '1';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when prepare_compute_4_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            if(reg_addition_subtraction_mode_q(0) = '0') then
                dsp2_b_en <= '0';
            else
                dsp2_b_en <= '1';
            end if;
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when compute_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '1';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            if(reg_addition_subtraction_mode_q(0) = '0') then
                dsp2_b_en <= '0';
            else
                dsp2_b_en <= '1';
            end if;
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_1_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '0';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            if(reg_addition_subtraction_mode_q(0) = '0') then
                dsp2_b_en <= '0';
            else
                dsp2_b_en <= '1';
            end if;
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_2_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '1';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '1';
            dsp1_a_rst <= '0';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '1';
            dsp1_c_rst <= '0';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            if(reg_addition_subtraction_mode_q(0) = '0') then
                dsp2_b_en <= '0';
            else
                dsp2_b_en <= '1';
            end if;
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_3_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '0';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '1';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            if(reg_addition_subtraction_mode_q(0) = '0') then
                dsp2_b_en <= '0';
            else
                dsp2_b_en <= '1';
            end if;
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_4_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            if(reg_addition_subtraction_mode_q(0) = '0') then
                dsp2_b_en <= '0';
            else
                dsp2_b_en <= '1';
            end if;
            dsp2_b_rst <= '1';
            dsp2_c_en <= '1';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_5_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '0';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '1';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '1';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when last_compute_6_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '1';
            reg_processor_free_d <= '1';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '0';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
        when finished_montgomery_addition_subtraction_no_reduction =>
            mem_write_enable_new_value <= '0';
            reg_processor_free_d <= '1';
            reg_addition_subtraction_mode_d <= "11";
            reg_addition_subtraction_mode_ce <= '0';
            reg_operands_size_ce <= '0';
            reg_variables_ce <= '0';
            counter_a_j_ce <= '0';
            counter_a_j_rst <= '1';
            counter_b_i_ce <= '0';
            counter_b_i_rst <= '1';
            address_n_ce <= '0';
            address_n_load <= '0';
            address_n_rst <= '1';
            address_new_p_ce <= '0';
            address_new_p_rst <= '1';
            dsp1_a_en <= '0';
            dsp1_a_rst <= '1';
            reg_b_ce <= '0';
            reg_b_rst <= '1';
            dsp1_c_en <= '0';
            dsp1_c_rst <= '1';
            dsp1_add_sub_mode <= '0';
            dsp1_reg_add_sub_mode_ce <= '0';
            dsp1_accumulation_mode <= '0';
            dsp1_reg_accumulation_mode_ce <= '0';
            dsp1_external_carry_in_mode <= '0';
            dsp1_reg_external_carry_in_mode_ce <= '0';
            dsp1_arshift_mode <= '0';
            dsp1_reg_arshift_mode_ce <= '0';
            dsp1_p_en <= '0';
            dsp1_p_rst <= '1';
            reg_m_ce <= '0';
            reg_m_rst <= '1';
            dsp2_b_en <= '0';
            dsp2_b_rst <= '1';
            dsp2_c_en <= '0';
            dsp2_c_rst <= '1';
            dsp2_add_sub_mode <= '0';
            dsp2_reg_add_sub_mode_ce <= '0';
            dsp2_accumulation_mode <= '0';
            dsp2_reg_accumulation_mode_ce <= '0';
            dsp2_external_carry_in_mode <= '0';
            dsp2_reg_external_carry_in_mode_ce <= '0';
            dsp2_arshift_mode <= '0';
            dsp2_reg_arshift_mode_ce <= '0';
            dsp2_p_en <= '0';
            dsp2_p_rst <= '1';
            sel_load_b_i <= '0';
            sel_value_m <= '0';
            sel_compare_counter_b_i <= '0';
    end case;
end process;


Update_Next_State : process (actual_state, start, instruction, counters_limit)
begin
    next_state <= reset;
    case (actual_state) is
        when reset =>
            next_state <= decode_instruction;
        when decode_instruction =>
            if(start = '1') then
                case (instruction) is
                    when "000" =>
                        next_state <= begin_montgomery_multiplication;
                    when "001" =>
                        next_state <= begin_montgomery_addition_subtraction_no_reduction;
                    when "010" =>
                        next_state <= begin_montgomery_addition_subtraction_no_reduction;
                    when "011" =>
                        next_state <= begin_montgomery_addition_subtraction_no_reduction;
                    when "111" =>
                        next_state <= decode_instruction;
                    when others =>
                        next_state <= decode_instruction;
                end case;
            else
                next_state <= decode_instruction;
            end if;
        when begin_montgomery_multiplication =>
            next_state <= begin_reset_counters_montgomery_multiplication;
        when begin_reset_counters_montgomery_multiplication =>
            next_state <= load_registers_1_first_iteration_montgomery_multiplication;
        when load_registers_1_first_iteration_montgomery_multiplication =>
            next_state <= load_registers_2_first_iteration_montgomery_multiplication;
        when load_registers_2_first_iteration_montgomery_multiplication =>
            next_state <= prepare_compute_m_1_first_iteration_montgomery_multiplication;
        when prepare_compute_m_1_first_iteration_montgomery_multiplication =>
            next_state <= prepare_compute_m_2_first_iteration_montgomery_multiplication;
        when prepare_compute_m_2_first_iteration_montgomery_multiplication =>
            next_state <= compute_m_first_iteration_montgomery_multiplication;
        when compute_m_first_iteration_montgomery_multiplication =>
            next_state <= prepare_compute_1_first_iteration_montgomery_multiplication;
        when prepare_compute_1_first_iteration_montgomery_multiplication =>
            next_state <= prepare_compute_2_first_iteration_montgomery_multiplication;
        when prepare_compute_2_first_iteration_montgomery_multiplication =>
            next_state <= prepare_compute_3_first_iteration_montgomery_multiplication;
        when prepare_compute_3_first_iteration_montgomery_multiplication =>
            next_state <= compute_first_iteration_montgomery_multiplication;
        when compute_first_iteration_montgomery_multiplication =>
            if(counters_limit = '1') then
                next_state <= last_compute_1_first_iteration_montgomery_multiplication;
            else
                next_state <= compute_first_iteration_montgomery_multiplication;
            end if;
        when last_compute_1_first_iteration_montgomery_multiplication =>
            next_state <= last_compute_2_first_iteration_montgomery_multiplication;
        when last_compute_2_first_iteration_montgomery_multiplication =>
            next_state <= last_compute_3_first_iteration_montgomery_multiplication;
        when last_compute_3_first_iteration_montgomery_multiplication =>
            next_state <= last_compute_4_remaining_iterations_montgomery_multiplication;
        when last_compute_4_remaining_iterations_montgomery_multiplication =>
            next_state <= prepare_compute_m_1_remaining_iterations_montgomery_multiplication;
        when prepare_compute_m_1_remaining_iterations_montgomery_multiplication =>
            next_state <= prepare_compute_m_2_remaining_iterations_montgomery_multiplication;
        when prepare_compute_m_2_remaining_iterations_montgomery_multiplication =>
            next_state <= compute_m_remaining_iterations_montgomery_multiplication;
        when compute_m_remaining_iterations_montgomery_multiplication =>
            next_state <= prepare_compute_1_remaining_iterations_montgomery_multiplication;
        when prepare_compute_1_remaining_iterations_montgomery_multiplication =>
            next_state <= prepare_compute_2_remaining_iterations_montgomery_multiplication;
        when prepare_compute_2_remaining_iterations_montgomery_multiplication =>
            next_state <= prepare_compute_3_remaining_iterations_montgomery_multiplication;
        when prepare_compute_3_remaining_iterations_montgomery_multiplication =>
            next_state <= compute_remaining_iterations_montgomery_multiplication;
        when compute_remaining_iterations_montgomery_multiplication =>
            if(counters_limit = '1') then
                next_state <= last_compute_1_remaining_iterations_montgomery_multiplication;
            else
                next_state <= compute_remaining_iterations_montgomery_multiplication;
            end if;
        when last_compute_1_remaining_iterations_montgomery_multiplication =>
            if(counters_limit = '1') then
                next_state <= last_compute_2_last_iterations_montgomery_multiplication;
            else
                next_state <= last_compute_2_remaining_iterations_montgomery_multiplication;
            end if;
        when last_compute_2_remaining_iterations_montgomery_multiplication =>
            next_state <= last_compute_3_remaining_iterations_montgomery_multiplication;
        when last_compute_3_remaining_iterations_montgomery_multiplication =>
            next_state <= last_compute_4_remaining_iterations_montgomery_multiplication;
        when last_compute_2_last_iterations_montgomery_multiplication =>
            next_state <= last_compute_3_last_iteration_montgomery_multiplication;
        when last_compute_3_last_iteration_montgomery_multiplication =>
            next_state <= last_compute_4_last_iteration_montgomery_multiplication;
        when last_compute_4_last_iteration_montgomery_multiplication =>
            next_state <= last_compute_5_last_iteration_montgomery_multiplication;
        when last_compute_5_last_iteration_montgomery_multiplication =>
            next_state <= last_compute_6_last_iteration_montgomery_multiplication;
        when last_compute_6_last_iteration_montgomery_multiplication =>
            next_state <= last_compute_7_last_iteration_montgomery_multiplication;
        when last_compute_7_last_iteration_montgomery_multiplication =>
            next_state <= finished_montgomery_multiplication;
        when finished_montgomery_multiplication =>
            next_state <= decode_instruction;
        when begin_montgomery_addition_subtraction_no_reduction =>
            next_state <= begin_reset_counters_montgomery_addition_subtraction_no_reduction;
        when begin_reset_counters_montgomery_addition_subtraction_no_reduction =>
            next_state <= prepare_compute_1_montgomery_addition_subtraction_no_reduction;
        when prepare_compute_1_montgomery_addition_subtraction_no_reduction =>
            next_state <= prepare_compute_2_montgomery_addition_subtraction_no_reduction;
        when prepare_compute_2_montgomery_addition_subtraction_no_reduction =>
            next_state <= prepare_compute_3_montgomery_addition_subtraction_no_reduction;
        when prepare_compute_3_montgomery_addition_subtraction_no_reduction =>
            next_state <= prepare_compute_4_montgomery_addition_subtraction_no_reduction;
        when prepare_compute_4_montgomery_addition_subtraction_no_reduction =>
            next_state <= compute_montgomery_addition_subtraction_no_reduction;
        when compute_montgomery_addition_subtraction_no_reduction =>
            if(counters_limit = '1') then
                next_state <= last_compute_1_montgomery_addition_subtraction_no_reduction;
            else
                next_state <= compute_montgomery_addition_subtraction_no_reduction;
            end if;
        when last_compute_1_montgomery_addition_subtraction_no_reduction =>
            next_state <= last_compute_2_montgomery_addition_subtraction_no_reduction;
        when last_compute_2_montgomery_addition_subtraction_no_reduction =>
            next_state <= last_compute_3_montgomery_addition_subtraction_no_reduction;
        when last_compute_3_montgomery_addition_subtraction_no_reduction =>
            next_state <= last_compute_4_montgomery_addition_subtraction_no_reduction;
        when last_compute_4_montgomery_addition_subtraction_no_reduction =>
            next_state <= last_compute_5_montgomery_addition_subtraction_no_reduction;
        when last_compute_5_montgomery_addition_subtraction_no_reduction =>
            next_state <= last_compute_6_montgomery_addition_subtraction_no_reduction;
        when last_compute_6_montgomery_addition_subtraction_no_reduction =>
            next_state <= finished_montgomery_addition_subtraction_no_reduction;
        when finished_montgomery_addition_subtraction_no_reduction =>
            next_state <= decode_instruction;
    end case;
end process;


reg_addition_subtraction_mode : register_rst_nbits
    Generic Map(
        size => 2
    )
    Port Map(
        d => reg_addition_subtraction_mode_d,
        clk => clk,
        ce => reg_addition_subtraction_mode_ce,
        rst => rst,
        rst_value => reg_addition_subtraction_mode_rst_value,
        q => reg_addition_subtraction_mode_q
    );

end Behavioral;